VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rdac3v_8bit
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rdac3v_8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 84.615 BY 156.255 ;
  PIN b0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 80.740 0.000 81.030 2.825 ;
    END
  END b0
  PIN b1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 72.600 0.000 72.890 2.825 ;
    END
  END b1
  PIN b2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 64.460 0.000 64.750 2.825 ;
    END
  END b2
  PIN b3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 56.320 0.000 56.610 2.825 ;
    END
  END b3
  PIN b4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 48.180 0.000 48.470 2.825 ;
    END
  END b4
  PIN b5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 40.040 0.000 40.330 2.825 ;
    END
  END b5
  PIN b6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 31.900 0.000 32.190 2.825 ;
    END
  END b6
  PIN b7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 23.760 0.000 24.050 2.825 ;
    END
  END b7
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.400000 ;
    ANTENNADIFFAREA 48.430000 ;
    PORT
      LAYER met2 ;
        RECT 34.360 153.635 35.635 156.255 ;
    END
  END out
  PIN vdd
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.005 0.000 3.105 156.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.495 31.695 84.615 33.000 ;
    END
  END vdd
  PIN vss
    ANTENNAGATEAREA 68.250000 ;
    ANTENNADIFFAREA 76.670097 ;
    PORT
      LAYER met3 ;
        RECT 82.225 124.185 84.175 127.715 ;
    END
    PORT
      LAYER met4 ;
	RECT 3.960 29.605 6.090 134.400 ;
        RECT 3.960 26.760 7.000 29.605 ;
        RECT 3.960 0.000 6.765 26.760 ;
        RECT 3.960 134.400 7.145 156.220 ;
    END
  END vss
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.702500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT 16.630 0.000 16.810 2.825 ;
    END
  END ena
  PIN dvdd
    ANTENNADIFFAREA 7.862400 ;
    PORT
      LAYER met2 ;
        RECT 11.810 0.000 13.535 2.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.120 0.000 78.030 7.250 ;
    END
  END dvdd
  PIN dvss
    ANTENNADIFFAREA 214.649200 ;
    PORT
      LAYER met2 ;
        RECT 9.155 0.000 11.050 8.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.705 0.000 84.615 7.270 ;
    END
  END dvss
  PIN Vhigh
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER met3 ;
        RECT 77.290 34.480 84.615 35.665 ;
    END
  END Vhigh
  PIN Vlow
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER met3 ;
        RECT 76.790 122.735 84.615 123.840 ;
    END
  END Vlow
  OBS
      LAYER nwell ;
        RECT 4.315 0.000 84.505 155.600 ;
      LAYER li1 ;
        RECT 4.545 0.330 84.075 156.215 ;
      LAYER met1 ;
        RECT 4.535 21.795 84.615 156.215 ;
        RECT 4.535 0.330 16.350 21.795 ;
        RECT 17.090 3.105 84.615 21.795 ;
        RECT 17.090 0.330 23.480 3.105 ;
        RECT 24.330 0.330 31.620 3.105 ;
        RECT 32.470 0.330 39.760 3.105 ;
        RECT 40.610 0.330 47.900 3.105 ;
        RECT 48.750 0.330 56.040 3.105 ;
        RECT 56.890 0.330 64.180 3.105 ;
        RECT 65.030 0.330 72.320 3.105 ;
        RECT 73.170 0.330 80.460 3.105 ;
        RECT 81.310 0.330 84.615 3.105 ;
      LAYER met2 ;
        RECT 0.000 153.355 34.080 155.980 ;
        RECT 35.915 153.355 84.615 155.980 ;
        RECT 0.000 8.350 84.615 153.355 ;
        RECT 0.000 0.610 8.875 8.350 ;
        RECT 11.330 3.265 84.615 8.350 ;
        RECT 11.330 0.610 11.530 3.265 ;
        RECT 13.815 0.610 84.615 3.265 ;
      LAYER met3 ;
        RECT 0.000 128.115 84.615 155.980 ;
        RECT 0.000 124.240 81.825 128.115 ;
        RECT 84.575 124.240 84.615 128.115 ;
        RECT 0.000 122.335 76.390 124.240 ;
        RECT 0.000 36.065 84.615 122.335 ;
        RECT 0.000 34.080 76.890 36.065 ;
        RECT 0.000 33.400 84.615 34.080 ;
        RECT 0.000 31.295 81.095 33.400 ;
        RECT 0.000 0.610 84.615 31.295 ;
      LAYER met4 ;
        RECT 7.575 134.000 84.615 138.710 ;
        RECT 7.165 27.270 84.615 134.000 ;
        RECT 7.165 7.670 84.615 27.270 ;
        RECT 7.165 7.650 82.305 7.670 ;
        RECT 7.165 7.250 75.720 7.650 ;
        RECT 78.430 7.250 82.305 7.650 ;
      LAYER met5 ;
        RECT 13.955 38.415 75.655 114.635 ;
  END
END sky130_ef_ip__rdac3v_8bit
END LIBRARY

