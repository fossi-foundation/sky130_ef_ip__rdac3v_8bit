magic
tech sky130A
magscale 1 2
timestamp 1740590524
<< dnwell >>
rect 1132 5855 16792 25830
<< nwell >>
rect 1023 25624 16901 25939
rect 1023 6061 1338 25624
rect 16586 6061 16901 25624
rect 1023 5746 16901 6061
<< pwell >>
rect 863 26224 16725 26558
<< mvpsubdiff >>
rect 909 26450 16687 26516
rect 909 26332 979 26450
rect 16595 26332 16687 26450
rect 909 26274 16687 26332
<< mvnsubdiff >>
rect 1089 25853 16835 25873
rect 1089 25819 1169 25853
rect 16755 25819 16835 25853
rect 1089 25799 16835 25819
rect 1089 25793 1163 25799
rect 1089 5892 1109 25793
rect 1143 5892 1163 25793
rect 1089 5886 1163 5892
rect 16761 25793 16835 25799
rect 16761 5892 16781 25793
rect 16815 5892 16835 25793
rect 16761 5886 16835 5892
rect 1089 5866 16835 5886
rect 1089 5832 1169 5866
rect 16755 5832 16835 5866
rect 1089 5812 16835 5832
<< mvpsubdiffcont >>
rect 979 26332 16595 26450
<< mvnsubdiffcont >>
rect 1169 25819 16755 25853
rect 1109 5892 1143 25793
rect 16781 5892 16815 25793
rect 1169 5832 16755 5866
<< locali >>
rect 909 26450 16687 26516
rect 909 26332 979 26450
rect 16595 26332 16687 26450
rect 909 26274 16687 26332
rect 1109 25819 1169 25853
rect 16755 25819 16815 25853
rect 1109 25793 1143 25819
rect 1109 5866 1143 5892
rect 16781 25793 16815 25819
rect 16781 5866 16815 5892
rect 1109 5832 1169 5866
rect 16755 5832 16815 5866
<< viali >>
rect 979 26332 16595 26450
rect 1181 25819 16745 25853
rect 1109 5903 1143 25782
rect 16781 5903 16815 25781
rect 1181 5832 16743 5866
<< metal1 >>
rect 16475 27048 16923 27050
rect 13577 27034 16923 27048
rect 13577 26972 16487 27034
rect 13559 26876 16487 26972
rect 16909 26876 16923 27034
rect 13559 26864 16923 26876
rect 13577 26862 16923 26864
rect 16751 26842 16923 26862
rect 16751 26514 16765 26842
rect 907 26450 16765 26514
rect 907 26332 979 26450
rect 16595 26332 16765 26450
rect 907 26290 16765 26332
rect 16911 26290 16923 26842
rect 907 26274 16923 26290
rect 1089 25853 16835 25873
rect 1089 25819 1181 25853
rect 16745 25819 16835 25853
rect 1089 25799 16835 25819
rect 1089 25782 1163 25799
rect 1089 5903 1109 25782
rect 1143 5903 1163 25782
rect 1250 25728 16696 25799
rect 16761 25781 16835 25799
rect 1250 25690 16692 25728
rect 1250 25544 1298 25690
rect 16664 25544 16692 25690
rect 1250 25504 16692 25544
rect 15440 25325 16064 25375
rect 15371 24469 15458 24475
rect 14971 24310 15371 24425
rect 15371 24260 15458 24266
rect 15371 7413 15458 7419
rect 14971 7254 15371 7369
rect 15371 7204 15458 7210
rect 15442 6304 16060 6354
rect 1242 6143 16684 6185
rect 1242 5997 1273 6143
rect 16639 5997 16684 6143
rect 1242 5957 16684 5997
rect 1089 5886 1163 5903
rect 16761 5903 16781 25781
rect 16815 5903 16835 25781
rect 16761 5886 16835 5903
rect 1089 5866 16835 5886
rect 1089 5832 1181 5866
rect 16743 5832 16835 5866
rect 1089 5812 16835 5832
rect 16106 5739 16314 5747
rect 15163 5661 15370 5669
rect 15162 5609 15163 5661
rect 13414 5585 13621 5597
rect 13413 5533 13414 5585
rect 11906 5433 12114 5445
rect 11905 5381 11906 5433
rect 10278 5281 10486 5291
rect 10277 5229 10278 5281
rect 8850 5129 9058 5142
rect 8850 5057 9058 5077
rect 7022 4977 7230 4986
rect 7021 4925 7022 4977
rect 6338 4825 6546 4835
rect 5394 4749 5602 4761
rect 5393 4697 5394 4749
rect 4710 4673 4918 4688
rect 3766 4597 3974 4610
rect 3765 4545 3766 4597
rect 3316 4523 3378 4533
rect 3766 4440 3974 4545
rect 4710 4440 4918 4621
rect 5394 4440 5602 4697
rect 6338 4440 6546 4773
rect 7022 4440 7230 4925
rect 7966 4901 8174 4913
rect 7966 4440 8174 4849
rect 8650 4770 9058 5057
rect 9594 5053 9802 5061
rect 8650 4440 8858 4770
rect 9594 4440 9802 5001
rect 10278 4440 10486 5229
rect 11222 5205 11430 5218
rect 11222 4440 11430 5153
rect 11906 4440 12114 5381
rect 12850 5357 13058 5370
rect 12850 4440 13058 5305
rect 13414 5335 13621 5533
rect 14478 5509 14686 5524
rect 13414 5108 13741 5335
rect 13534 4440 13741 5108
rect 14478 4440 14686 5457
rect 15163 4446 15370 5609
rect 16106 4440 16314 5687
rect 3316 4293 3378 4303
rect 1831 1792 2460 1812
rect 1831 1614 1853 1792
rect 2441 1614 2460 1792
rect 1831 1593 2460 1614
rect 3326 244 3362 4293
rect 3234 238 3442 244
rect 3234 184 3246 238
rect 3430 184 3442 238
rect 3234 178 3442 184
rect 4698 236 4906 242
rect 4698 182 4710 236
rect 4894 182 4906 236
rect 4698 176 4906 182
rect 6326 236 6534 242
rect 6326 182 6338 236
rect 6522 182 6534 236
rect 6326 176 6534 182
rect 7954 236 8162 242
rect 7954 182 7966 236
rect 8150 182 8162 236
rect 7954 176 8162 182
rect 9582 236 9790 242
rect 9582 182 9594 236
rect 9778 182 9790 236
rect 9582 176 9790 182
rect 11210 236 11418 242
rect 11210 182 11222 236
rect 11406 182 11418 236
rect 11210 176 11418 182
rect 12838 236 13046 242
rect 12838 182 12850 236
rect 13034 182 13046 236
rect 12838 176 13046 182
rect 14466 236 14674 242
rect 14466 182 14478 236
rect 14662 182 14674 236
rect 14466 176 14674 182
rect 16094 236 16302 242
rect 16094 182 16106 236
rect 16290 182 16302 236
rect 16094 176 16302 182
rect 4752 67 4810 176
rect 6380 67 6438 176
rect 8008 67 8066 176
rect 9636 67 9694 176
rect 11264 67 11322 176
rect 12892 67 12950 176
rect 14520 67 14578 176
rect 16148 67 16206 176
<< via1 >>
rect 16487 26876 16909 27034
rect 16765 26290 16911 26842
rect 1298 25544 16664 25690
rect 15371 24266 15458 24469
rect 15371 7210 15458 7413
rect 1273 5997 16639 6143
rect 16106 5687 16314 5739
rect 15163 5609 15370 5661
rect 13414 5533 13621 5585
rect 11906 5381 12114 5433
rect 10278 5229 10486 5281
rect 8850 5077 9058 5129
rect 7022 4925 7230 4977
rect 6338 4773 6546 4825
rect 5394 4697 5602 4749
rect 4710 4621 4918 4673
rect 3766 4545 3974 4597
rect 3316 4303 3378 4523
rect 7966 4849 8174 4901
rect 9594 5001 9802 5053
rect 11222 5153 11430 5205
rect 12850 5305 13058 5357
rect 14478 5457 14686 5509
rect 1853 1614 2441 1792
rect 3246 184 3430 238
rect 4710 182 4894 236
rect 6338 182 6522 236
rect 7966 182 8150 236
rect 9594 182 9778 236
rect 11222 182 11406 236
rect 12850 182 13034 236
rect 14478 182 14662 236
rect 16106 182 16290 236
<< metal2 >>
rect 6872 30997 7127 31251
rect 13845 31192 16189 31196
rect 13845 31134 16827 31192
rect 13845 27436 16497 31134
rect 16775 27436 16827 31134
rect 13845 27386 16827 27436
rect 3793 26800 3833 27136
rect 4281 26894 4299 27136
rect 4787 26894 4799 27136
rect 4281 26866 4799 26894
rect 665 26760 3833 26800
rect 0 25705 625 25734
rect 0 25182 23 25705
rect 607 25182 625 25705
rect 0 25148 625 25182
rect 11 21395 595 21414
rect 11 15815 18 21395
rect 578 15815 595 21395
rect 11 15791 593 15815
rect 533 15016 593 15791
rect 533 14960 535 15016
rect 591 14960 593 15016
rect 533 14958 593 14960
rect 535 14951 591 14958
rect 7 14824 538 14843
rect 7 12434 24 14824
rect 514 12434 538 14824
rect 7 12407 538 12434
rect 665 4513 701 26760
rect 1427 26062 1613 26068
rect 1427 26000 1439 26062
rect 1601 26050 1613 26062
rect 5597 26050 5641 27138
rect 13845 26132 16189 27386
rect 16475 27034 16923 27050
rect 16475 26876 16487 27034
rect 16909 26876 16923 27034
rect 16475 26862 16923 26876
rect 16751 26842 16923 26862
rect 16751 26290 16765 26842
rect 16911 26290 16923 26842
rect 1601 26006 5641 26050
rect 1601 26000 1613 26006
rect 1427 25994 1613 26000
rect 1249 25718 16692 25732
rect 1249 25714 12873 25718
rect 1249 25690 1765 25714
rect 2097 25712 12873 25714
rect 2097 25690 2323 25712
rect 2559 25708 12873 25712
rect 2559 25690 5929 25708
rect 6165 25690 12873 25708
rect 13283 25690 16692 25718
rect 1249 25544 1298 25690
rect 16664 25544 16692 25690
rect 1249 25538 1765 25544
rect 2097 25538 2323 25544
rect 1249 25534 2323 25538
rect 2559 25534 5929 25544
rect 1249 25530 5929 25534
rect 6165 25532 12873 25544
rect 13283 25532 16692 25544
rect 6165 25530 16692 25532
rect 1249 25504 16692 25530
rect 1250 25422 1538 25504
rect 2820 25428 3045 25504
rect 4327 25431 4552 25504
rect 5834 25428 6059 25504
rect 7341 25429 7566 25504
rect 8848 25431 9073 25504
rect 10355 25427 10580 25504
rect 11862 25428 12087 25504
rect 13369 25429 13594 25504
rect 14876 25428 15101 25504
rect 16383 25431 16684 25504
rect 746 4589 782 19417
rect 822 4665 858 19297
rect 898 4741 934 21552
rect 974 4817 1010 21431
rect 1250 6248 1401 25422
rect 15271 24693 15358 24702
rect 15358 24552 15458 24589
rect 15271 24502 15458 24552
rect 15371 24469 15458 24502
rect 15371 24260 15458 24266
rect 3348 23653 3404 23736
rect 3348 15125 3404 15207
rect 15371 7413 15458 7419
rect 15371 7087 15458 7210
rect 15371 6937 15458 6946
rect 16521 6800 16684 25431
rect 16671 6600 16684 6800
rect 2070 6185 2295 6249
rect 3577 6185 3802 6249
rect 5084 6185 5309 6252
rect 6591 6185 6816 6252
rect 8098 6185 8323 6250
rect 9605 6185 9830 6250
rect 11112 6185 11337 6255
rect 12619 6185 12844 6250
rect 14126 6185 14351 6257
rect 15633 6185 15858 6259
rect 16521 6248 16684 6600
rect 1242 6162 16684 6185
rect 1242 5977 1267 6162
rect 2762 6143 16684 6162
rect 16639 5997 16684 6143
rect 2762 5977 16684 5997
rect 1242 5957 16684 5977
rect 16099 5731 16106 5739
rect 16014 5729 16106 5731
rect 2923 5695 16106 5729
rect 2923 5693 16045 5695
rect 16099 5687 16106 5695
rect 16314 5731 16320 5739
rect 16314 5695 16329 5731
rect 16314 5687 16320 5695
rect 15155 5653 15163 5661
rect 2923 5617 15163 5653
rect 15155 5609 15163 5617
rect 15370 5609 15376 5661
rect 13406 5577 13414 5585
rect 2923 5541 13414 5577
rect 13406 5533 13414 5541
rect 13621 5577 13627 5585
rect 13621 5541 13762 5577
rect 13621 5533 13627 5541
rect 14471 5501 14478 5509
rect 2923 5465 14478 5501
rect 14471 5457 14478 5465
rect 14686 5501 14692 5509
rect 14686 5465 14701 5501
rect 14686 5457 14692 5465
rect 11898 5425 11906 5433
rect 2923 5389 11906 5425
rect 11898 5381 11906 5389
rect 12114 5425 12120 5433
rect 12114 5389 12257 5425
rect 12114 5381 12120 5389
rect 12843 5349 12850 5357
rect 2923 5313 12850 5349
rect 12843 5305 12850 5313
rect 13058 5349 13064 5357
rect 13058 5313 13071 5349
rect 13058 5305 13064 5313
rect 10270 5273 10278 5281
rect 2923 5237 10278 5273
rect 10270 5229 10278 5237
rect 10486 5273 10492 5281
rect 10486 5237 10501 5273
rect 10486 5229 10492 5237
rect 11215 5197 11222 5205
rect 2923 5161 11222 5197
rect 11215 5153 11222 5161
rect 11430 5197 11436 5205
rect 11430 5161 11443 5197
rect 11430 5153 11436 5161
rect 8842 5121 8850 5129
rect 2923 5085 8850 5121
rect 8842 5077 8850 5085
rect 9058 5121 9064 5129
rect 9058 5085 14793 5121
rect 9058 5077 9064 5085
rect 9587 5045 9594 5053
rect 2923 5009 9594 5045
rect 9587 5001 9594 5009
rect 9802 5045 9808 5053
rect 9802 5009 14534 5045
rect 9802 5001 9808 5009
rect 7014 4969 7022 4977
rect 2923 4933 7022 4969
rect 7014 4925 7022 4933
rect 7230 4969 7236 4977
rect 7230 4933 7239 4969
rect 7230 4925 7236 4933
rect 7959 4893 7966 4901
rect 2923 4857 7966 4893
rect 7959 4849 7966 4857
rect 8174 4893 8180 4901
rect 8174 4857 8191 4893
rect 8174 4849 8180 4857
rect 6331 4817 6338 4825
rect 974 4781 6338 4817
rect 6331 4773 6338 4781
rect 6546 4817 6552 4825
rect 6546 4781 6561 4817
rect 6546 4773 6552 4781
rect 5386 4741 5394 4749
rect 898 4705 5394 4741
rect 5386 4697 5394 4705
rect 5602 4741 5608 4749
rect 5602 4705 5619 4741
rect 5602 4697 5608 4705
rect 4704 4665 4710 4673
rect 822 4629 4710 4665
rect 4704 4621 4710 4629
rect 4918 4665 4925 4673
rect 4918 4629 4940 4665
rect 4918 4621 4925 4629
rect 3758 4589 3766 4597
rect 746 4553 3766 4589
rect 3758 4545 3766 4553
rect 3974 4589 3980 4597
rect 3974 4553 3985 4589
rect 3974 4545 3980 4553
rect 3306 4513 3316 4523
rect 665 4477 3316 4513
rect 3306 4303 3316 4477
rect 3378 4303 3388 4523
rect 2574 4007 3491 4022
rect 2574 3652 2601 4007
rect 3250 3652 3491 4007
rect 2574 3643 3491 3652
rect 16751 1811 16923 26290
rect 1831 1792 16923 1811
rect 1831 1614 1853 1792
rect 2441 1784 16923 1792
rect 2441 1614 16576 1784
rect 1831 1454 16576 1614
rect 16886 1454 16923 1784
rect 1831 1432 16923 1454
rect 1831 0 2210 1432
rect 2574 1210 3494 1222
rect 2574 855 2601 1210
rect 3250 855 3494 1210
rect 2574 843 3494 855
rect 15224 597 15606 598
rect 2362 568 16894 597
rect 2362 304 15248 568
rect 2362 0 2707 304
rect 3234 238 3442 244
rect 3234 184 3246 238
rect 3430 184 3442 238
rect 3234 178 3442 184
rect 4698 236 4906 242
rect 4698 182 4710 236
rect 4894 182 4906 236
rect 3326 0 3362 178
rect 4698 176 4906 182
rect 6326 236 6534 242
rect 6326 182 6338 236
rect 6522 182 6534 236
rect 6326 176 6534 182
rect 7954 236 8162 242
rect 7954 182 7966 236
rect 8150 182 8162 236
rect 7954 176 8162 182
rect 9582 236 9790 242
rect 9582 182 9594 236
rect 9778 182 9790 236
rect 9582 176 9790 182
rect 11210 236 11418 242
rect 11210 182 11222 236
rect 11406 182 11418 236
rect 11210 176 11418 182
rect 12838 236 13046 242
rect 12838 182 12850 236
rect 13034 182 13046 236
rect 12838 176 13046 182
rect 14466 236 14674 242
rect 14466 182 14478 236
rect 14662 182 14674 236
rect 14466 176 14674 182
rect 4752 0 4810 176
rect 6380 0 6438 176
rect 8008 0 8066 176
rect 9636 0 9694 176
rect 11264 0 11322 176
rect 12892 0 12950 176
rect 14520 0 14578 176
rect 15224 150 15248 304
rect 15572 304 16894 568
rect 15572 150 15606 304
rect 16094 236 16302 242
rect 16094 182 16106 236
rect 16290 182 16302 236
rect 16094 176 16302 182
rect 15224 122 15606 150
rect 16148 0 16206 176
<< via2 >>
rect 16497 27436 16775 31134
rect 4299 26894 4787 27346
rect 23 25182 607 25705
rect 18 15815 578 21395
rect 535 14960 591 15016
rect 24 12434 514 14824
rect 1439 26000 1601 26062
rect 5941 27134 13253 27306
rect 1765 25690 2097 25714
rect 2323 25690 2559 25712
rect 5929 25690 6165 25708
rect 12873 25690 13283 25718
rect 1765 25544 2097 25690
rect 2323 25544 2559 25690
rect 5929 25544 6165 25690
rect 12873 25544 13283 25690
rect 1765 25538 2097 25544
rect 2323 25534 2559 25544
rect 5929 25530 6165 25544
rect 12873 25532 13283 25544
rect 15640 24846 15851 25031
rect 15271 24552 15358 24693
rect 15371 6946 15458 7087
rect 16514 6600 16671 6800
rect 1267 6143 2762 6162
rect 1267 5997 1273 6143
rect 1273 5997 2762 6143
rect 1267 5977 2762 5997
rect 2601 3652 3250 4007
rect 16576 1454 16886 1784
rect 2601 855 3250 1210
rect 15248 150 15572 568
<< metal3 >>
rect 1 27742 621 27786
rect 1 26178 43 27742
rect 579 26698 621 27742
rect 4271 27346 4815 27366
rect 4271 26894 4299 27346
rect 4787 26894 4815 27346
rect 4271 26868 4815 26894
rect 5913 27306 13297 27340
rect 5913 27134 5941 27306
rect 13253 27134 13297 27306
rect 5913 26698 13297 27134
rect 579 26688 13297 26698
rect 13845 27266 16187 31196
rect 16447 31134 16827 31192
rect 16447 27436 16497 31134
rect 16775 28234 16827 31134
rect 16775 27436 16829 28234
rect 16447 27386 16829 27436
rect 13845 26688 16189 27266
rect 579 26666 16189 26688
rect 579 26178 1515 26666
rect 1 26164 1515 26178
rect 2529 26638 16189 26666
rect 2529 26168 5963 26638
rect 13235 26168 16189 26638
rect 2529 26164 16189 26168
rect 1 26136 16189 26164
rect 1487 26134 2117 26136
rect 1427 26062 1613 26068
rect 1427 26000 1439 26062
rect 1601 26000 1613 26062
rect 1427 25994 1613 26000
rect 0 25705 639 25734
rect 0 25182 23 25705
rect 607 25182 639 25705
rect 1429 25444 1497 25994
rect 1749 25714 2117 26134
rect 1749 25538 1765 25714
rect 2097 25538 2117 25714
rect 1749 25516 2117 25538
rect 2305 25712 2573 26136
rect 2305 25534 2323 25712
rect 2559 25534 2573 25712
rect 2305 25516 2573 25534
rect 5913 25708 6181 26136
rect 5913 25530 5929 25708
rect 6165 25530 6181 25708
rect 5913 25516 6181 25530
rect 12861 25718 13299 26136
rect 13845 26132 16189 26136
rect 16449 25874 16829 27386
rect 12861 25532 12873 25718
rect 13283 25532 13299 25718
rect 12861 25516 13299 25532
rect 16445 25865 16835 25874
rect 16445 25543 16454 25865
rect 16826 25543 16835 25865
rect 0 25148 639 25182
rect 1 23546 639 25148
rect 1419 25426 1509 25444
rect 1419 25160 1431 25426
rect 1497 25160 1509 25426
rect 1419 25140 1509 25160
rect 16445 25197 16835 25543
rect 16445 25039 16923 25197
rect 15633 25031 16923 25039
rect 15633 24846 15640 25031
rect 15851 24846 16923 25031
rect 15633 24837 16923 24846
rect 15266 24693 16923 24768
rect 15266 24552 15271 24693
rect 15358 24552 16923 24693
rect 15266 24547 16923 24552
rect 845 23744 1195 23754
rect 1195 23622 1333 23672
rect 845 23612 1333 23622
rect 1 23486 1337 23546
rect 1 23389 639 23486
rect 1 21395 53 23389
rect 1 15815 18 21395
rect 586 15860 639 23389
rect 3198 22412 3283 22474
rect 3223 22351 3283 22412
rect 3072 22010 3132 22291
rect 3223 22285 3446 22351
rect 3072 21950 3392 22010
rect 2300 21611 2869 21671
rect 884 21480 1337 21540
rect 956 21354 1337 21414
rect 1501 19790 3566 19850
rect 2300 19479 2868 19539
rect 730 19348 1337 19408
rect 802 19222 1337 19282
rect 3198 18148 3283 18210
rect 3223 18087 3283 18148
rect 3072 17746 3132 18027
rect 3223 18021 3446 18087
rect 3072 17686 3392 17746
rect 2300 17347 2869 17407
rect 958 17216 1337 17276
rect 880 17090 1337 17150
rect 578 15815 639 15860
rect 1 15791 639 15815
rect 1197 15520 1529 15580
rect 223 15084 1355 15144
rect 223 14857 283 15084
rect 530 15018 596 15021
rect 530 15016 1355 15018
rect 530 14960 535 15016
rect 591 14960 1355 15016
rect 530 14958 1355 14960
rect 530 14955 596 14958
rect 10 14824 535 14857
rect 10 12434 24 14824
rect 514 12434 535 14824
rect 3198 13884 3283 13946
rect 3223 13823 3283 13884
rect 3072 13482 3132 13763
rect 3223 13757 3446 13823
rect 3072 13422 3392 13482
rect 2300 13083 2869 13143
rect 883 12952 1355 13012
rect 955 12826 1355 12886
rect 10 6194 535 12434
rect 1510 11262 3575 11322
rect 2300 10951 2868 11011
rect 807 10820 1355 10880
rect 724 10694 1355 10754
rect 3204 9620 3283 9682
rect 3223 9559 3283 9620
rect 3072 9218 3132 9495
rect 3223 9493 3367 9559
rect 3072 9158 3307 9218
rect 2301 8819 2871 8879
rect 957 8688 1355 8748
rect 877 8562 1355 8622
rect 15366 7087 16923 7133
rect 15366 6946 15371 7087
rect 15458 6946 16923 7087
rect 15366 6896 16923 6946
rect 16258 6800 16923 6814
rect 16258 6600 16514 6800
rect 16671 6600 16923 6800
rect 16258 6587 16923 6600
rect 16299 6339 16923 6587
rect 10 6170 2788 6194
rect 3136 6192 3196 6195
rect 3265 6192 3325 6195
rect 3394 6192 3454 6195
rect 3523 6192 3583 6195
rect 3790 6192 3850 6195
rect 3919 6192 3979 6195
rect 4048 6192 4108 6195
rect 4177 6192 4237 6195
rect 4643 6192 4703 6195
rect 4772 6192 4832 6195
rect 4901 6192 4961 6195
rect 5030 6192 5090 6195
rect 5297 6192 5357 6195
rect 5426 6192 5486 6195
rect 5555 6192 5615 6195
rect 5684 6192 5744 6195
rect 6150 6192 6210 6195
rect 6279 6192 6339 6195
rect 6408 6192 6468 6195
rect 6537 6192 6597 6195
rect 6804 6192 6864 6195
rect 6933 6192 6993 6195
rect 7062 6192 7122 6195
rect 7191 6192 7251 6195
rect 7657 6192 7717 6195
rect 7786 6192 7846 6195
rect 7915 6192 7975 6195
rect 8044 6192 8104 6195
rect 8311 6192 8371 6195
rect 8440 6192 8500 6195
rect 8569 6192 8629 6195
rect 8698 6192 8758 6195
rect 9164 6192 9224 6195
rect 9293 6192 9353 6195
rect 9422 6192 9482 6195
rect 9551 6192 9611 6195
rect 9818 6192 9878 6195
rect 9947 6192 10007 6195
rect 10076 6192 10136 6195
rect 10205 6192 10265 6195
rect 10671 6192 10731 6195
rect 10800 6192 10860 6195
rect 10929 6192 10989 6195
rect 11058 6192 11118 6195
rect 11325 6192 11385 6195
rect 11454 6192 11514 6195
rect 11583 6192 11643 6195
rect 11712 6192 11772 6195
rect 12178 6192 12238 6195
rect 12307 6192 12367 6195
rect 12436 6192 12496 6195
rect 12565 6192 12625 6195
rect 12832 6192 12892 6195
rect 12961 6192 13021 6195
rect 13090 6192 13150 6195
rect 13219 6192 13279 6195
rect 13685 6192 13745 6195
rect 13814 6192 13874 6195
rect 13943 6192 14003 6195
rect 14072 6192 14132 6195
rect 14339 6192 14399 6195
rect 14468 6192 14528 6195
rect 14597 6192 14657 6195
rect 14726 6192 14786 6195
rect 10 5374 811 6170
rect 1202 6162 2788 6170
rect 1202 5977 1267 6162
rect 2762 5977 2788 6162
rect 1202 5948 2788 5977
rect 3134 6186 3198 6192
rect 1202 5886 1648 5948
rect 3134 5942 3198 5948
rect 3263 6186 3327 6192
rect 3263 5942 3327 5948
rect 3392 6186 3456 6192
rect 3392 5942 3456 5948
rect 3521 6186 3585 6192
rect 3521 5942 3585 5948
rect 3788 6186 3852 6192
rect 3788 5942 3852 5948
rect 3917 6186 3981 6192
rect 3917 5942 3981 5948
rect 4046 6186 4110 6192
rect 4046 5942 4110 5948
rect 4175 6186 4239 6192
rect 4175 5942 4239 5948
rect 4641 6186 4705 6192
rect 4641 5942 4705 5948
rect 4770 6186 4834 6192
rect 4770 5942 4834 5948
rect 4899 6186 4963 6192
rect 4899 5942 4963 5948
rect 5028 6186 5092 6192
rect 5028 5942 5092 5948
rect 5295 6186 5359 6192
rect 5295 5942 5359 5948
rect 5424 6186 5488 6192
rect 5424 5942 5488 5948
rect 5553 6186 5617 6192
rect 5553 5942 5617 5948
rect 5682 6186 5746 6192
rect 5682 5942 5746 5948
rect 6148 6186 6212 6192
rect 6148 5942 6212 5948
rect 6277 6186 6341 6192
rect 6277 5942 6341 5948
rect 6406 6186 6470 6192
rect 6406 5942 6470 5948
rect 6535 6186 6599 6192
rect 6535 5942 6599 5948
rect 6802 6186 6866 6192
rect 6802 5942 6866 5948
rect 6931 6186 6995 6192
rect 6931 5942 6995 5948
rect 7060 6186 7124 6192
rect 7060 5942 7124 5948
rect 7189 6186 7253 6192
rect 7189 5942 7253 5948
rect 7655 6186 7719 6192
rect 7655 5942 7719 5948
rect 7784 6186 7848 6192
rect 7784 5942 7848 5948
rect 7913 6186 7977 6192
rect 7913 5942 7977 5948
rect 8042 6186 8106 6192
rect 8042 5942 8106 5948
rect 8309 6186 8373 6192
rect 8309 5942 8373 5948
rect 8438 6186 8502 6192
rect 8438 5942 8502 5948
rect 8567 6186 8631 6192
rect 8567 5942 8631 5948
rect 8696 6186 8760 6192
rect 8696 5942 8760 5948
rect 9162 6186 9226 6192
rect 9162 5942 9226 5948
rect 9291 6186 9355 6192
rect 9291 5942 9355 5948
rect 9420 6186 9484 6192
rect 9420 5942 9484 5948
rect 9549 6186 9613 6192
rect 9549 5942 9613 5948
rect 9816 6186 9880 6192
rect 9816 5942 9880 5948
rect 9945 6186 10009 6192
rect 9945 5942 10009 5948
rect 10074 6186 10138 6192
rect 10074 5942 10138 5948
rect 10203 6186 10267 6192
rect 10203 5942 10267 5948
rect 10669 6186 10733 6192
rect 10669 5942 10733 5948
rect 10798 6186 10862 6192
rect 10798 5942 10862 5948
rect 10927 6186 10991 6192
rect 10927 5942 10991 5948
rect 11056 6186 11120 6192
rect 11056 5942 11120 5948
rect 11323 6186 11387 6192
rect 11323 5942 11387 5948
rect 11452 6186 11516 6192
rect 11452 5942 11516 5948
rect 11581 6186 11645 6192
rect 11581 5942 11645 5948
rect 11710 6186 11774 6192
rect 11710 5942 11774 5948
rect 12176 6186 12240 6192
rect 12176 5942 12240 5948
rect 12305 6186 12369 6192
rect 12305 5942 12369 5948
rect 12434 6186 12498 6192
rect 12434 5942 12498 5948
rect 12563 6186 12627 6192
rect 12563 5942 12627 5948
rect 12830 6186 12894 6192
rect 12830 5942 12894 5948
rect 12959 6186 13023 6192
rect 12959 5942 13023 5948
rect 13088 6186 13152 6192
rect 13088 5942 13152 5948
rect 13217 6186 13281 6192
rect 13217 5942 13281 5948
rect 13683 6186 13747 6192
rect 13683 5942 13747 5948
rect 13812 6186 13876 6192
rect 13812 5942 13876 5948
rect 13941 6186 14005 6192
rect 13941 5942 14005 5948
rect 14070 6186 14134 6192
rect 14070 5942 14134 5948
rect 14337 6186 14401 6192
rect 14337 5942 14401 5948
rect 14466 6186 14530 6192
rect 14466 5942 14530 5948
rect 14595 6186 14659 6192
rect 14595 5942 14659 5948
rect 14724 6186 14788 6192
rect 14724 5942 14788 5948
rect 1202 5388 1323 5886
rect 1613 5388 1648 5886
rect 1202 5374 1648 5388
rect 10 5352 1648 5374
rect 3136 4916 3196 5942
rect 3265 5595 3325 5942
rect 3394 4911 3454 5942
rect 3523 5671 3583 5942
rect 3790 5593 3850 5942
rect 3919 5440 3979 5942
rect 4048 5670 4108 5942
rect 4177 5521 4237 5942
rect 4643 5444 4703 5942
rect 4772 5667 4832 5942
rect 4901 5518 4961 5942
rect 5030 5595 5090 5942
rect 5297 5671 5357 5942
rect 5426 5294 5486 5942
rect 5555 5597 5615 5942
rect 5684 5367 5744 5942
rect 6150 5287 6210 5942
rect 6279 5594 6339 5942
rect 6408 5369 6468 5942
rect 6537 5670 6597 5942
rect 6804 5594 6864 5942
rect 6933 5517 6993 5942
rect 7062 5670 7122 5942
rect 7191 5446 7251 5942
rect 7657 5517 7717 5942
rect 7786 5670 7846 5942
rect 7915 5443 7975 5942
rect 8044 5594 8104 5942
rect 8311 5668 8371 5942
rect 8440 5212 8500 5942
rect 8569 5594 8629 5942
rect 8698 5142 8758 5942
rect 9164 5213 9224 5942
rect 9293 5594 9353 5942
rect 9422 5139 9482 5942
rect 9551 5665 9611 5942
rect 9818 5593 9878 5942
rect 9947 5441 10007 5942
rect 10076 5671 10136 5942
rect 10205 5517 10265 5942
rect 10671 5444 10731 5942
rect 10800 5671 10860 5942
rect 10929 5516 10989 5942
rect 11058 5591 11118 5942
rect 11325 5671 11385 5942
rect 11454 5370 11514 5942
rect 11583 5594 11643 5942
rect 11712 5293 11772 5942
rect 12178 5367 12238 5942
rect 12307 5595 12367 5942
rect 12436 5292 12496 5942
rect 12565 5668 12625 5942
rect 12832 5595 12892 5942
rect 12961 5525 13021 5942
rect 13090 5671 13150 5942
rect 13219 5443 13279 5942
rect 13685 5524 13745 5942
rect 13814 5674 13874 5942
rect 13943 5439 14003 5942
rect 14072 5597 14132 5942
rect 14339 5665 14399 5942
rect 14468 5066 14528 5942
rect 14597 5598 14657 5942
rect 14726 5068 14786 5942
rect 16299 5855 16719 6339
rect 16299 5523 16309 5855
rect 16713 5523 16719 5855
rect 16299 5516 16719 5523
rect 1895 4323 2537 4324
rect 1 4309 3261 4323
rect 1 4302 1914 4309
rect 1 3658 17 4302
rect 597 3658 1914 4302
rect 1 3655 1914 3658
rect 2505 4007 3261 4309
rect 2505 3655 2601 4007
rect 1 3652 2601 3655
rect 3250 3652 3261 4007
rect 1 3639 3261 3652
rect 2593 1210 3261 3639
rect 2593 855 2601 1210
rect 3250 855 3261 1210
rect 2593 826 3261 855
rect 15224 1794 15606 1826
rect 15224 1450 15246 1794
rect 15578 1450 15606 1794
rect 15224 568 15606 1450
rect 16540 1784 16922 1810
rect 16540 1454 16576 1784
rect 16886 1454 16922 1784
rect 16540 1432 16922 1454
rect 15224 150 15248 568
rect 15572 150 15606 568
rect 15224 122 15606 150
<< via3 >>
rect 43 26178 579 27742
rect 4299 26894 4787 27346
rect 1515 26164 2529 26666
rect 5963 26168 13235 26638
rect 16454 25543 16826 25865
rect 1431 25160 1497 25426
rect 845 23622 1195 23744
rect 53 21395 586 23389
rect 53 15860 578 21395
rect 578 15860 586 21395
rect 811 5374 1202 6170
rect 3134 5948 3198 6186
rect 3263 5948 3327 6186
rect 3392 5948 3456 6186
rect 3521 5948 3585 6186
rect 3788 5948 3852 6186
rect 3917 5948 3981 6186
rect 4046 5948 4110 6186
rect 4175 5948 4239 6186
rect 4641 5948 4705 6186
rect 4770 5948 4834 6186
rect 4899 5948 4963 6186
rect 5028 5948 5092 6186
rect 5295 5948 5359 6186
rect 5424 5948 5488 6186
rect 5553 5948 5617 6186
rect 5682 5948 5746 6186
rect 6148 5948 6212 6186
rect 6277 5948 6341 6186
rect 6406 5948 6470 6186
rect 6535 5948 6599 6186
rect 6802 5948 6866 6186
rect 6931 5948 6995 6186
rect 7060 5948 7124 6186
rect 7189 5948 7253 6186
rect 7655 5948 7719 6186
rect 7784 5948 7848 6186
rect 7913 5948 7977 6186
rect 8042 5948 8106 6186
rect 8309 5948 8373 6186
rect 8438 5948 8502 6186
rect 8567 5948 8631 6186
rect 8696 5948 8760 6186
rect 9162 5948 9226 6186
rect 9291 5948 9355 6186
rect 9420 5948 9484 6186
rect 9549 5948 9613 6186
rect 9816 5948 9880 6186
rect 9945 5948 10009 6186
rect 10074 5948 10138 6186
rect 10203 5948 10267 6186
rect 10669 5948 10733 6186
rect 10798 5948 10862 6186
rect 10927 5948 10991 6186
rect 11056 5948 11120 6186
rect 11323 5948 11387 6186
rect 11452 5948 11516 6186
rect 11581 5948 11645 6186
rect 11710 5948 11774 6186
rect 12176 5948 12240 6186
rect 12305 5948 12369 6186
rect 12434 5948 12498 6186
rect 12563 5948 12627 6186
rect 12830 5948 12894 6186
rect 12959 5948 13023 6186
rect 13088 5948 13152 6186
rect 13217 5948 13281 6186
rect 13683 5948 13747 6186
rect 13812 5948 13876 6186
rect 13941 5948 14005 6186
rect 14070 5948 14134 6186
rect 14337 5948 14401 6186
rect 14466 5948 14530 6186
rect 14595 5948 14659 6186
rect 14724 5948 14788 6186
rect 1323 5388 1613 5886
rect 16309 5523 16713 5855
rect 17 3658 597 4302
rect 1914 3655 2505 4309
rect 15246 1450 15578 1794
rect 16576 1454 16886 1784
<< metal4 >>
rect 1 27742 621 31244
rect 1 26178 43 27742
rect 579 26178 621 27742
rect 1 23389 621 26178
rect 1 15860 53 23389
rect 586 15860 621 23389
rect 1 4302 621 15860
rect 1 3658 17 4302
rect 597 3658 621 4302
rect 1 0 621 3658
rect 792 27362 1429 31244
rect 792 27346 4809 27362
rect 792 26894 4299 27346
rect 4787 26894 4809 27346
rect 792 26880 4809 26894
rect 792 25875 1218 26880
rect 1485 26666 13299 26692
rect 1485 26164 1515 26666
rect 2529 26638 13299 26666
rect 2529 26168 5963 26638
rect 13235 26168 13299 26638
rect 2529 26164 13299 26168
rect 1485 26136 13299 26164
rect 792 25865 16835 25875
rect 792 25543 16454 25865
rect 16826 25543 16835 25865
rect 792 25534 16835 25543
rect 792 23744 1218 25534
rect 1419 25426 1510 25444
rect 1419 25160 1431 25426
rect 1497 25160 1510 25426
rect 1419 25140 1510 25160
rect 792 23622 845 23744
rect 1195 23622 1218 23744
rect 792 6170 1218 23622
rect 1450 11261 1510 25140
rect 2156 17484 2216 21527
rect 3649 20535 3709 22527
rect 3649 19313 3709 19700
rect 3649 16268 3709 18260
rect 2156 8962 2216 13005
rect 3649 12001 3709 13993
rect 3649 10785 3709 11172
rect 3649 7741 3709 9733
rect 3139 7290 3195 7385
rect 3396 7291 3452 7386
rect 3136 6187 3196 6255
rect 3265 6187 3325 6255
rect 3394 6187 3454 6255
rect 3523 6187 3583 6255
rect 3790 6187 3850 6255
rect 3919 6187 3979 6255
rect 4048 6187 4108 6255
rect 4177 6187 4237 6255
rect 4643 6187 4703 6255
rect 4772 6187 4832 6255
rect 4901 6187 4961 6255
rect 5030 6187 5090 6255
rect 5297 6187 5357 6255
rect 5426 6187 5486 6255
rect 5555 6187 5615 6255
rect 5684 6187 5744 6255
rect 6150 6187 6210 6255
rect 6279 6187 6339 6255
rect 6408 6187 6468 6255
rect 6537 6187 6597 6255
rect 6804 6187 6864 6255
rect 6933 6187 6993 6255
rect 7062 6187 7122 6255
rect 7191 6187 7251 6255
rect 7657 6187 7717 6255
rect 7786 6187 7846 6255
rect 7915 6187 7975 6255
rect 8044 6187 8104 6255
rect 8311 6187 8371 6255
rect 8440 6187 8500 6255
rect 8569 6187 8629 6255
rect 8698 6187 8758 6255
rect 9164 6187 9224 6255
rect 9293 6187 9353 6255
rect 9422 6187 9482 6255
rect 9551 6187 9611 6255
rect 9818 6187 9878 6255
rect 9947 6187 10007 6255
rect 10076 6187 10136 6255
rect 10205 6187 10265 6255
rect 10671 6187 10731 6255
rect 10800 6187 10860 6255
rect 10929 6187 10989 6255
rect 11058 6187 11118 6255
rect 11325 6187 11385 6255
rect 11454 6187 11514 6255
rect 11583 6187 11643 6255
rect 11712 6187 11772 6255
rect 12178 6187 12238 6255
rect 12307 6187 12367 6255
rect 12436 6187 12496 6255
rect 12565 6187 12625 6255
rect 12832 6187 12892 6255
rect 12961 6187 13021 6255
rect 13090 6187 13150 6255
rect 13219 6187 13279 6255
rect 13685 6187 13745 6255
rect 13814 6187 13874 6255
rect 13943 6187 14003 6255
rect 14072 6187 14132 6255
rect 14339 6187 14399 6255
rect 14468 6187 14528 6255
rect 14597 6187 14657 6255
rect 14726 6187 14786 6255
rect 792 5374 811 6170
rect 1202 5921 1218 6170
rect 3133 6186 3199 6187
rect 3133 5948 3134 6186
rect 3198 5948 3199 6186
rect 3133 5947 3199 5948
rect 3262 6186 3328 6187
rect 3262 5948 3263 6186
rect 3327 5948 3328 6186
rect 3262 5947 3328 5948
rect 3391 6186 3457 6187
rect 3391 5948 3392 6186
rect 3456 5948 3457 6186
rect 3391 5947 3457 5948
rect 3520 6186 3586 6187
rect 3520 5948 3521 6186
rect 3585 5948 3586 6186
rect 3520 5947 3586 5948
rect 3787 6186 3853 6187
rect 3787 5948 3788 6186
rect 3852 5948 3853 6186
rect 3787 5947 3853 5948
rect 3916 6186 3982 6187
rect 3916 5948 3917 6186
rect 3981 5948 3982 6186
rect 3916 5947 3982 5948
rect 4045 6186 4111 6187
rect 4045 5948 4046 6186
rect 4110 5948 4111 6186
rect 4045 5947 4111 5948
rect 4174 6186 4240 6187
rect 4174 5948 4175 6186
rect 4239 5948 4240 6186
rect 4174 5947 4240 5948
rect 4640 6186 4706 6187
rect 4640 5948 4641 6186
rect 4705 5948 4706 6186
rect 4640 5947 4706 5948
rect 4769 6186 4835 6187
rect 4769 5948 4770 6186
rect 4834 5948 4835 6186
rect 4769 5947 4835 5948
rect 4898 6186 4964 6187
rect 4898 5948 4899 6186
rect 4963 5948 4964 6186
rect 4898 5947 4964 5948
rect 5027 6186 5093 6187
rect 5027 5948 5028 6186
rect 5092 5948 5093 6186
rect 5027 5947 5093 5948
rect 5294 6186 5360 6187
rect 5294 5948 5295 6186
rect 5359 5948 5360 6186
rect 5294 5947 5360 5948
rect 5423 6186 5489 6187
rect 5423 5948 5424 6186
rect 5488 5948 5489 6186
rect 5423 5947 5489 5948
rect 5552 6186 5618 6187
rect 5552 5948 5553 6186
rect 5617 5948 5618 6186
rect 5552 5947 5618 5948
rect 5681 6186 5747 6187
rect 5681 5948 5682 6186
rect 5746 5948 5747 6186
rect 5681 5947 5747 5948
rect 6147 6186 6213 6187
rect 6147 5948 6148 6186
rect 6212 5948 6213 6186
rect 6147 5947 6213 5948
rect 6276 6186 6342 6187
rect 6276 5948 6277 6186
rect 6341 5948 6342 6186
rect 6276 5947 6342 5948
rect 6405 6186 6471 6187
rect 6405 5948 6406 6186
rect 6470 5948 6471 6186
rect 6405 5947 6471 5948
rect 6534 6186 6600 6187
rect 6534 5948 6535 6186
rect 6599 5948 6600 6186
rect 6534 5947 6600 5948
rect 6801 6186 6867 6187
rect 6801 5948 6802 6186
rect 6866 5948 6867 6186
rect 6801 5947 6867 5948
rect 6930 6186 6996 6187
rect 6930 5948 6931 6186
rect 6995 5948 6996 6186
rect 6930 5947 6996 5948
rect 7059 6186 7125 6187
rect 7059 5948 7060 6186
rect 7124 5948 7125 6186
rect 7059 5947 7125 5948
rect 7188 6186 7254 6187
rect 7188 5948 7189 6186
rect 7253 5948 7254 6186
rect 7188 5947 7254 5948
rect 7654 6186 7720 6187
rect 7654 5948 7655 6186
rect 7719 5948 7720 6186
rect 7654 5947 7720 5948
rect 7783 6186 7849 6187
rect 7783 5948 7784 6186
rect 7848 5948 7849 6186
rect 7783 5947 7849 5948
rect 7912 6186 7978 6187
rect 7912 5948 7913 6186
rect 7977 5948 7978 6186
rect 7912 5947 7978 5948
rect 8041 6186 8107 6187
rect 8041 5948 8042 6186
rect 8106 5948 8107 6186
rect 8041 5947 8107 5948
rect 8308 6186 8374 6187
rect 8308 5948 8309 6186
rect 8373 5948 8374 6186
rect 8308 5947 8374 5948
rect 8437 6186 8503 6187
rect 8437 5948 8438 6186
rect 8502 5948 8503 6186
rect 8437 5947 8503 5948
rect 8566 6186 8632 6187
rect 8566 5948 8567 6186
rect 8631 5948 8632 6186
rect 8566 5947 8632 5948
rect 8695 6186 8761 6187
rect 8695 5948 8696 6186
rect 8760 5948 8761 6186
rect 8695 5947 8761 5948
rect 9161 6186 9227 6187
rect 9161 5948 9162 6186
rect 9226 5948 9227 6186
rect 9161 5947 9227 5948
rect 9290 6186 9356 6187
rect 9290 5948 9291 6186
rect 9355 5948 9356 6186
rect 9290 5947 9356 5948
rect 9419 6186 9485 6187
rect 9419 5948 9420 6186
rect 9484 5948 9485 6186
rect 9419 5947 9485 5948
rect 9548 6186 9614 6187
rect 9548 5948 9549 6186
rect 9613 5948 9614 6186
rect 9548 5947 9614 5948
rect 9815 6186 9881 6187
rect 9815 5948 9816 6186
rect 9880 5948 9881 6186
rect 9815 5947 9881 5948
rect 9944 6186 10010 6187
rect 9944 5948 9945 6186
rect 10009 5948 10010 6186
rect 9944 5947 10010 5948
rect 10073 6186 10139 6187
rect 10073 5948 10074 6186
rect 10138 5948 10139 6186
rect 10073 5947 10139 5948
rect 10202 6186 10268 6187
rect 10202 5948 10203 6186
rect 10267 5948 10268 6186
rect 10202 5947 10268 5948
rect 10668 6186 10734 6187
rect 10668 5948 10669 6186
rect 10733 5948 10734 6186
rect 10668 5947 10734 5948
rect 10797 6186 10863 6187
rect 10797 5948 10798 6186
rect 10862 5948 10863 6186
rect 10797 5947 10863 5948
rect 10926 6186 10992 6187
rect 10926 5948 10927 6186
rect 10991 5948 10992 6186
rect 10926 5947 10992 5948
rect 11055 6186 11121 6187
rect 11055 5948 11056 6186
rect 11120 5948 11121 6186
rect 11055 5947 11121 5948
rect 11322 6186 11388 6187
rect 11322 5948 11323 6186
rect 11387 5948 11388 6186
rect 11322 5947 11388 5948
rect 11451 6186 11517 6187
rect 11451 5948 11452 6186
rect 11516 5948 11517 6186
rect 11451 5947 11517 5948
rect 11580 6186 11646 6187
rect 11580 5948 11581 6186
rect 11645 5948 11646 6186
rect 11580 5947 11646 5948
rect 11709 6186 11775 6187
rect 11709 5948 11710 6186
rect 11774 5948 11775 6186
rect 11709 5947 11775 5948
rect 12175 6186 12241 6187
rect 12175 5948 12176 6186
rect 12240 5948 12241 6186
rect 12175 5947 12241 5948
rect 12304 6186 12370 6187
rect 12304 5948 12305 6186
rect 12369 5948 12370 6186
rect 12304 5947 12370 5948
rect 12433 6186 12499 6187
rect 12433 5948 12434 6186
rect 12498 5948 12499 6186
rect 12433 5947 12499 5948
rect 12562 6186 12628 6187
rect 12562 5948 12563 6186
rect 12627 5948 12628 6186
rect 12562 5947 12628 5948
rect 12829 6186 12895 6187
rect 12829 5948 12830 6186
rect 12894 5948 12895 6186
rect 12829 5947 12895 5948
rect 12958 6186 13024 6187
rect 12958 5948 12959 6186
rect 13023 5948 13024 6186
rect 12958 5947 13024 5948
rect 13087 6186 13153 6187
rect 13087 5948 13088 6186
rect 13152 5948 13153 6186
rect 13087 5947 13153 5948
rect 13216 6186 13282 6187
rect 13216 5948 13217 6186
rect 13281 5948 13282 6186
rect 13216 5947 13282 5948
rect 13682 6186 13748 6187
rect 13682 5948 13683 6186
rect 13747 5948 13748 6186
rect 13682 5947 13748 5948
rect 13811 6186 13877 6187
rect 13811 5948 13812 6186
rect 13876 5948 13877 6186
rect 13811 5947 13877 5948
rect 13940 6186 14006 6187
rect 13940 5948 13941 6186
rect 14005 5948 14006 6186
rect 13940 5947 14006 5948
rect 14069 6186 14135 6187
rect 14069 5948 14070 6186
rect 14134 5948 14135 6186
rect 14069 5947 14135 5948
rect 14336 6186 14402 6187
rect 14336 5948 14337 6186
rect 14401 5948 14402 6186
rect 14336 5947 14402 5948
rect 14465 6186 14531 6187
rect 14465 5948 14466 6186
rect 14530 5948 14531 6186
rect 14465 5947 14531 5948
rect 14594 6186 14660 6187
rect 14594 5948 14595 6186
rect 14659 5948 14660 6186
rect 14594 5947 14660 5948
rect 14723 6186 14789 6187
rect 14723 5948 14724 6186
rect 14788 5948 14789 6186
rect 14723 5947 14789 5948
rect 3136 5941 3196 5947
rect 3265 5941 3325 5947
rect 3394 5941 3454 5947
rect 3523 5941 3583 5947
rect 3790 5941 3850 5947
rect 3919 5941 3979 5947
rect 4048 5941 4108 5947
rect 4177 5941 4237 5947
rect 4643 5941 4703 5947
rect 4772 5941 4832 5947
rect 4901 5941 4961 5947
rect 5030 5941 5090 5947
rect 5297 5941 5357 5947
rect 5426 5941 5486 5947
rect 5555 5941 5615 5947
rect 5684 5941 5744 5947
rect 6150 5941 6210 5947
rect 6279 5941 6339 5947
rect 6408 5941 6468 5947
rect 6537 5941 6597 5947
rect 6804 5941 6864 5947
rect 6933 5941 6993 5947
rect 7062 5941 7122 5947
rect 7191 5941 7251 5947
rect 7657 5941 7717 5947
rect 7786 5941 7846 5947
rect 7915 5941 7975 5947
rect 8044 5941 8104 5947
rect 8311 5941 8371 5947
rect 8440 5941 8500 5947
rect 8569 5941 8629 5947
rect 8698 5941 8758 5947
rect 9164 5941 9224 5947
rect 9293 5941 9353 5947
rect 9422 5941 9482 5947
rect 9551 5941 9611 5947
rect 9818 5941 9878 5947
rect 9947 5941 10007 5947
rect 10076 5941 10136 5947
rect 10205 5941 10265 5947
rect 10671 5941 10731 5947
rect 10800 5941 10860 5947
rect 10929 5941 10989 5947
rect 11058 5941 11118 5947
rect 11325 5941 11385 5947
rect 11454 5941 11514 5947
rect 11583 5941 11643 5947
rect 11712 5941 11772 5947
rect 12178 5941 12238 5947
rect 12307 5941 12367 5947
rect 12436 5941 12496 5947
rect 12565 5941 12625 5947
rect 12832 5941 12892 5947
rect 12961 5941 13021 5947
rect 13090 5941 13150 5947
rect 13219 5941 13279 5947
rect 13685 5941 13745 5947
rect 13814 5941 13874 5947
rect 13943 5941 14003 5947
rect 14072 5941 14132 5947
rect 14339 5941 14399 5947
rect 14468 5941 14528 5947
rect 14597 5941 14657 5947
rect 14726 5941 14786 5947
rect 1202 5886 1648 5921
rect 1202 5388 1323 5886
rect 1613 5388 1648 5886
rect 1202 5374 1648 5388
rect 792 5352 1648 5374
rect 1901 5855 16835 5869
rect 1901 5523 16309 5855
rect 16713 5523 16835 5855
rect 1901 5517 16835 5523
rect 792 0 1353 5352
rect 1901 4309 2521 5517
rect 1901 3655 1914 4309
rect 2505 3655 2521 4309
rect 1901 3632 2521 3655
rect 15224 1794 15606 4429
rect 15224 1450 15246 1794
rect 15578 1450 15606 1794
rect 15224 0 15606 1450
rect 16541 1784 16923 4429
rect 16541 1454 16576 1784
rect 16886 1454 16923 1784
rect 16541 0 16923 1454
use dac_3v_column  dac_3v_column_0
timestamp 1653060931
transform 0 -1 16579 1 0 7331
box -20 -7 1049 15264
use dac_3v_column  dac_3v_column_1
timestamp 1653060931
transform 0 -1 16579 1 0 9463
box -20 -7 1049 15264
use dac_3v_column  dac_3v_column_2
timestamp 1653060931
transform 0 -1 16579 1 0 11595
box -20 -7 1049 15264
use dac_3v_column  dac_3v_column_3
timestamp 1653060931
transform 0 -1 16579 1 0 13727
box -20 -7 1049 15264
use dac_3v_column  dac_3v_column_4
timestamp 1653060931
transform 0 -1 16579 1 0 15859
box -20 -7 1049 15264
use dac_3v_column  dac_3v_column_5
timestamp 1653060931
transform 0 -1 16579 1 0 17991
box -20 -7 1049 15264
use dac_3v_column  dac_3v_column_6
timestamp 1653060931
transform 0 -1 16579 1 0 20123
box -20 -7 1049 15264
use dac_3v_column  dac_3v_column_7
timestamp 1653060931
transform 0 -1 16579 1 0 22255
box -20 -7 1049 15264
use dac_3v_column_dummy  dac_3v_column_dummy_0
timestamp 1653061945
transform 0 -1 16579 1 0 6266
box -18 -7 1049 15272
use dac_3v_column_dummy  dac_3v_column_dummy_1
timestamp 1653061945
transform 0 -1 16579 1 0 24386
box -18 -7 1049 15272
use dac_3v_column_odd  dac_3v_column_odd_0
timestamp 1653060931
transform 0 -1 16579 1 0 8398
box -20 -7 1049 15263
use dac_3v_column_odd  dac_3v_column_odd_1
timestamp 1653060931
transform 0 -1 16579 1 0 10530
box -20 -7 1049 15263
use dac_3v_column_odd  dac_3v_column_odd_2
timestamp 1653060931
transform 0 -1 16579 1 0 12662
box -20 -7 1049 15263
use dac_3v_column_odd  dac_3v_column_odd_3
timestamp 1653060931
transform 0 -1 16579 1 0 14794
box -20 -7 1049 15263
use dac_3v_column_odd  dac_3v_column_odd_4
timestamp 1653060931
transform 0 -1 16579 1 0 16926
box -20 -7 1049 15263
use dac_3v_column_odd  dac_3v_column_odd_5
timestamp 1653060931
transform 0 -1 16579 1 0 19058
box -20 -7 1049 15263
use dac_3v_column_odd  dac_3v_column_odd_6
timestamp 1653060931
transform 0 -1 16579 1 0 21190
box -20 -7 1049 15263
use dac_3v_column_odd  dac_3v_column_odd_7
timestamp 1653060931
transform 0 -1 16579 1 0 23322
box -20 -7 1049 15263
use follower_amp  follower_amp_0 ../ip/sky130_ef_ip__samplehold/mag
timestamp 1740434940
transform 0 1 2540 1 0 26866
box 0 -1436 4377 11129
use level_shifter_array  level_shifter_array_0
timestamp 1652995732
transform 0 -1 16589 1 0 23
box -23 -10 4908 13105
use m2m3contact  m2m3contact_0
timestamp 1652924542
transform 1 0 14443 0 1 4224
box 276 844 350 997
use m2m3contact  m2m3contact_1
timestamp 1652924542
transform 1 0 14315 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_2
timestamp 1652924542
transform 1 0 14056 0 1 4831
box 276 844 350 997
use m2m3contact  m2m3contact_3
timestamp 1652924542
transform 1 0 13402 0 1 4679
box 276 844 350 997
use m2m3contact  m2m3contact_4
timestamp 1652924542
transform 1 0 13660 0 1 4604
box 276 844 350 997
use m2m3contact  m2m3contact_5
timestamp 1652924542
transform 1 0 12807 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_6
timestamp 1652924542
transform 1 0 12548 0 1 4755
box 276 844 350 997
use m2m3contact  m2m3contact_7
timestamp 1652924542
transform 1 0 11300 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_8
timestamp 1652924542
transform 1 0 11041 0 1 4831
box 276 844 350 997
use m2m3contact  m2m3contact_9
timestamp 1652924542
transform 1 0 12153 0 1 4452
box 276 844 350 997
use m2m3contact  m2m3contact_10
timestamp 1652924542
transform 1 0 11895 0 1 4527
box 276 844 350 997
use m2m3contact  m2m3contact_11
timestamp 1652924542
transform 1 0 8286 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_12
timestamp 1652924542
transform 1 0 8027 0 1 4831
box 276 844 350 997
use m2m3contact  m2m3contact_13
timestamp 1652924542
transform 1 0 5272 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_14
timestamp 1652924542
transform 1 0 5013 0 1 4831
box 276 844 350 997
use m2m3contact  m2m3contact_15
timestamp 1652924542
transform 1 0 9534 0 1 4755
box 276 844 350 997
use m2m3contact  m2m3contact_16
timestamp 1652924542
transform 1 0 9793 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_17
timestamp 1652924542
transform 1 0 6520 0 1 4755
box 276 844 350 997
use m2m3contact  m2m3contact_18
timestamp 1652924542
transform 1 0 6779 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_19
timestamp 1652924542
transform 1 0 3506 0 1 4755
box 276 844 350 997
use m2m3contact  m2m3contact_20
timestamp 1652924542
transform 1 0 3765 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_21
timestamp 1652924542
transform 1 0 10646 0 1 4680
box 276 844 350 997
use m2m3contact  m2m3contact_22
timestamp 1652924542
transform 1 0 10388 0 1 4603
box 276 844 350 997
use m2m3contact  m2m3contact_23
timestamp 1652924542
transform 1 0 9139 0 1 4300
box 276 844 350 997
use m2m3contact  m2m3contact_24
timestamp 1652924542
transform 1 0 8881 0 1 4375
box 276 844 350 997
use m2m3contact  m2m3contact_25
timestamp 1652924542
transform 1 0 7632 0 1 4604
box 276 844 350 997
use m2m3contact  m2m3contact_26
timestamp 1652924542
transform 1 0 7374 0 1 4679
box 276 844 350 997
use m2m3contact  m2m3contact_27
timestamp 1652924542
transform 1 0 6125 0 1 4528
box 276 844 350 997
use m2m3contact  m2m3contact_28
timestamp 1652924542
transform 1 0 5867 0 1 4451
box 276 844 350 997
use m2m3contact  m2m3contact_29
timestamp 1652924542
transform 1 0 4618 0 1 4680
box 276 844 350 997
use m2m3contact  m2m3contact_30
timestamp 1652924542
transform 1 0 4360 0 1 4603
box 276 844 350 997
use m2m3contact  m2m3contact_31
timestamp 1652924542
transform 1 0 3111 0 1 3996
box 276 844 350 997
use m2m3contact  m2m3contact_32
timestamp 1652924542
transform 1 0 2853 0 1 4071
box 276 844 350 997
use m2m3contact  m2m3contact_33
timestamp 1652924542
transform 1 0 14185 0 1 4148
box 276 844 350 997
use m2m3contact  m2m3contact_34
timestamp 1652924542
transform 1 0 13789 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_35
timestamp 1652924542
transform 1 0 13531 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_36
timestamp 1652924542
transform 1 0 12282 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_37
timestamp 1652924542
transform 1 0 12024 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_38
timestamp 1652924542
transform 1 0 9268 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_39
timestamp 1652924542
transform 1 0 9010 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_40
timestamp 1652924542
transform 1 0 6254 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_41
timestamp 1652924542
transform 1 0 5996 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_42
timestamp 1652924542
transform 1 0 3240 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_43
timestamp 1652924542
transform 1 0 2982 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_44
timestamp 1652924542
transform 1 0 10775 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_45
timestamp 1652924542
transform 1 0 10517 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_46
timestamp 1652924542
transform 1 0 7761 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_47
timestamp 1652924542
transform 1 0 7503 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_48
timestamp 1652924542
transform 1 0 4747 0 1 4756
box 276 844 350 997
use m2m3contact  m2m3contact_49
timestamp 1652924542
transform 1 0 4489 0 1 4832
box 276 844 350 997
use m2m3contact  m2m3contact_50
timestamp 1652924542
transform 1 0 12936 0 1 4604
box 276 844 350 997
use m2m3contact  m2m3contact_51
timestamp 1652924542
transform 1 0 12678 0 1 4680
box 276 844 350 997
use m2m3contact  m2m3contact_52
timestamp 1652924542
transform 1 0 11429 0 1 4452
box 276 844 350 997
use m2m3contact  m2m3contact_53
timestamp 1652924542
transform 1 0 11171 0 1 4528
box 276 844 350 997
use m2m3contact  m2m3contact_54
timestamp 1652924542
transform 1 0 9922 0 1 4680
box 276 844 350 997
use m2m3contact  m2m3contact_55
timestamp 1652924542
transform 1 0 9664 0 1 4604
box 276 844 350 997
use m2m3contact  m2m3contact_56
timestamp 1652924542
transform 1 0 8415 0 1 4300
box 276 844 350 997
use m2m3contact  m2m3contact_57
timestamp 1652924542
transform 1 0 8157 0 1 4376
box 276 844 350 997
use m2m3contact  m2m3contact_58
timestamp 1652924542
transform 1 0 6908 0 1 4604
box 276 844 350 997
use m2m3contact  m2m3contact_59
timestamp 1652924542
transform 1 0 6650 0 1 4680
box 276 844 350 997
use m2m3contact  m2m3contact_60
timestamp 1652924542
transform 1 0 5401 0 1 4528
box 276 844 350 997
use m2m3contact  m2m3contact_61
timestamp 1652924542
transform 1 0 5143 0 1 4452
box 276 844 350 997
use m2m3contact  m2m3contact_62
timestamp 1652924542
transform 1 0 3636 0 1 4604
box 276 844 350 997
use m2m3contact  m2m3contact_63
timestamp 1652924542
transform 1 0 3894 0 1 4680
box 276 844 350 997
use m2m3contact  m2m3contact_64
timestamp 1652924542
transform 0 -1 1873 1 0 8405
box 276 844 350 997
use m2m3contact  m2m3contact_65
timestamp 1652924542
transform 0 -1 1795 1 0 8279
box 276 844 350 997
use m2m3contact  m2m3contact_66
timestamp 1652924542
transform 0 -1 1643 1 0 10411
box 276 844 350 997
use m2m3contact  m2m3contact_67
timestamp 1652924542
transform 0 -1 1721 1 0 10537
box 276 844 350 997
use m2m3contact  m2m3contact_68
timestamp 1652924542
transform 0 -1 1871 1 0 12543
box 276 844 350 997
use m2m3contact  m2m3contact_69
timestamp 1652924542
transform 0 -1 1797 1 0 12669
box 276 844 350 997
use m2m3contact  m2m3contact_72
timestamp 1652924542
transform 0 -1 1795 1 0 16807
box 276 844 350 997
use m2m3contact  m2m3contact_73
timestamp 1652924542
transform 0 -1 1873 1 0 16933
box 276 844 350 997
use m2m3contact  m2m3contact_74
timestamp 1652924542
transform 0 -1 1719 1 0 18939
box 276 844 350 997
use m2m3contact  m2m3contact_75
timestamp 1652924542
transform 0 1 -116 1 0 19065
box 276 844 350 997
use m2m3contact  m2m3contact_76
timestamp 1652924542
transform 0 -1 1871 1 0 21071
box 276 844 350 997
use m2m3contact  m2m3contact_77
timestamp 1652924542
transform 0 -1 1797 1 0 21197
box 276 844 350 997
use m3m4contact  m3m4contact_0
timestamp 1652924542
transform 0 -1 10662 -1 0 7257
box -258 7458 -104 7613
use m3m4contact  m3m4contact_1
timestamp 1652924542
transform 0 -1 10920 -1 0 7257
box -258 7458 -104 7613
use m3m4contact  m3m4contact_2
timestamp 1652924542
transform 0 -1 10662 -1 0 11521
box -258 7458 -104 7613
use m3m4contact  m3m4contact_3
timestamp 1652924542
transform 0 -1 10920 -1 0 11521
box -258 7458 -104 7613
use m3m4contact  m3m4contact_4
timestamp 1652924542
transform 0 -1 10662 -1 0 15785
box -258 7458 -104 7613
use m3m4contact  m3m4contact_5
timestamp 1652924542
transform 0 -1 10920 -1 0 15785
box -258 7458 -104 7613
use m3m4contact  m3m4contact_6
timestamp 1652924542
transform 0 -1 10662 -1 0 20049
box -258 7458 -104 7613
use m3m4contact  m3m4contact_7
timestamp 1652924542
transform 0 -1 10920 -1 0 20049
box -258 7458 -104 7613
use m3m4contact  m3m4contact_8
timestamp 1652924542
transform 0 1 -4330 1 0 9789
box -258 7458 -104 7613
use m3m4contact  m3m4contact_9
timestamp 1652924542
transform 0 -1 10920 1 0 9325
box -258 7458 -104 7613
use m3m4contact  m3m4contact_10
timestamp 1652924542
transform 0 -1 10920 1 0 13589
box -258 7458 -104 7613
use m3m4contact  m3m4contact_11
timestamp 1652924542
transform 0 1 -4330 1 0 14053
box -258 7458 -104 7613
use m3m4contact  m3m4contact_12
timestamp 1652924542
transform 0 -1 10920 1 0 17853
box -258 7458 -104 7613
use m3m4contact  m3m4contact_13
timestamp 1652924542
transform 0 1 -4330 1 0 18317
box -258 7458 -104 7613
use m3m4contact  m3m4contact_14
timestamp 1652924542
transform 0 -1 10920 1 0 22117
box -258 7458 -104 7613
use m3m4contact  m3m4contact_15
timestamp 1652924542
transform 0 1 -4330 1 0 22581
box -258 7458 -104 7613
use m3m4contact  m3m4contact_16
timestamp 1652924542
transform 0 1 -5310 -1 0 8712
box -258 7458 -104 7613
use m3m4contact  m3m4contact_17
timestamp 1652924542
transform 0 1 -5310 1 0 13250
box -258 7458 -104 7613
use m3m4contact  m3m4contact_18
timestamp 1652924542
transform 0 1 -5310 -1 0 17240
box -258 7458 -104 7613
use m3m4contact  m3m4contact_19
timestamp 1652924542
transform 0 1 -5310 1 0 21778
box -258 7458 -104 7613
use m3m4contact  m3m4contact_20
timestamp 1652924542
transform 0 1 -5310 1 0 11118
box -258 7458 -104 7613
use m3m4contact  m3m4contact_21
timestamp 1652924542
transform 0 1 -5310 1 0 19646
box -258 7458 -104 7613
use m3m4contact  m3m4contact_22
timestamp 1652924542
transform 0 -1 11175 1 0 11429
box -258 7458 -104 7613
use m3m4contact  m3m4contact_23
timestamp 1652924542
transform 0 -1 11175 1 0 19957
box -258 7458 -104 7613
use m3m4contact  m3m4contact_24
timestamp 1652924542
transform 0 1 -6016 -1 0 11155
box -258 7458 -104 7613
use m3m4contact  m3m4contact_25
timestamp 1652924542
transform 0 1 -6016 -1 0 15413
box -258 7458 -104 7613
use m3m4contact  m3m4contact_26
timestamp 1652924542
transform 0 1 -6016 1 0 19957
box -258 7458 -104 7613
use m3m4contact  m3m4contact_27
timestamp 1652924542
transform 0 -1 11175 1 0 15687
box -258 7458 -104 7613
<< labels >>
flabel metal2 16148 0 16206 182 0 FreeSans 400 90 0 0 b[0]
port 1 nsew signal input
flabel metal2 14520 0 14578 182 0 FreeSans 400 270 0 0 b[1]
port 2 nsew signal input
flabel metal2 12892 0 12950 182 0 FreeSans 400 270 0 0 b[2]
port 3 nsew signal input
flabel metal2 11264 0 11322 182 0 FreeSans 400 270 0 0 b[3]
port 4 nsew signal input
flabel metal2 9636 0 9694 182 0 FreeSans 400 270 0 0 b[4]
port 5 nsew signal input
flabel metal2 8008 0 8066 182 0 FreeSans 400 270 0 0 b[5]
port 6 nsew signal input
flabel metal2 6380 0 6438 182 0 FreeSans 400 270 0 0 b[6]
port 7 nsew signal input
flabel metal2 4752 0 4810 182 0 FreeSans 400 270 0 0 b[7]
port 8 nsew signal input
flabel metal2 3326 0 3362 184 0 FreeSans 320 270 0 0 ena
port 12 nsew signal input
flabel metal4 s 1 0 621 31244 0 FreeSans 1600 270 0 0 avdd
port 10 nsew power bidirectional
flabel metal2 1831 0 2210 1614 0 FreeSans 1600 270 0 0 dvss
port 14 nsew ground bidirectional
flabel metal2 2362 0 2707 597 0 FreeSans 1600 270 0 0 dvdd
port 13 nsew power bidirectional
flabel metal3 15458 6896 16923 7133 0 FreeSans 480 270 0 0 Vhigh
port 15 nsew analog bidirectional
flabel metal3 s 16299 6339 16923 6814 0 FreeSans 400 270 0 0 avdd
port 10 nsew power bidirectional
flabel metal3 15358 24547 16923 24768 0 FreeSans 480 90 0 0 Vlow
port 16 nsew analog bidirectional
flabel metal3 16445 24837 16923 25197 0 FreeSans 400 270 0 0 avss
port 11 nsew ground bidirectional
flabel metal4 3169 7332 3169 7332 0 FreeSans 240 270 0 0 b5a
flabel metal4 3424 7332 3424 7332 0 FreeSans 240 270 0 0 b5b
flabel metal3 1263 15545 1263 15545 0 FreeSans 240 0 0 0 out_unbuf
flabel metal2 3005 4570 3005 4570 0 FreeSans 400 0 0 0 b7b
flabel metal2 3009 4722 3009 4722 0 FreeSans 400 0 0 0 b6b
flabel metal2 3008 4875 3008 4875 0 FreeSans 400 0 0 0 b5b
flabel metal2 3006 5024 3006 5024 0 FreeSans 400 0 0 0 b4b
flabel metal2 3003 5179 3003 5179 0 FreeSans 400 0 0 0 b3b
flabel metal2 3004 5328 3004 5328 0 FreeSans 400 0 0 0 b2b
flabel metal2 3016 5483 3016 5483 0 FreeSans 400 0 0 0 b1b
flabel metal2 3004 5634 3004 5634 0 FreeSans 400 0 0 0 b0b
flabel metal2 3004 4647 3004 4647 0 FreeSans 400 0 0 0 b7a
flabel metal2 3005 4799 3005 4799 0 FreeSans 400 0 0 0 b6a
flabel metal2 3009 4952 3009 4952 0 FreeSans 400 0 0 0 b5a
flabel metal2 3007 5103 3007 5103 0 FreeSans 400 0 0 0 b4a
flabel metal2 3005 5256 3005 5256 0 FreeSans 400 0 0 0 b3a
flabel metal2 3004 5406 3004 5406 0 FreeSans 400 0 0 0 b2a
flabel metal2 3016 5560 3016 5560 0 FreeSans 400 0 0 0 b1a
flabel metal2 3009 5711 3009 5711 0 FreeSans 400 0 0 0 b0a
flabel metal3 1267 8596 1267 8596 0 FreeSans 240 90 0 0 b6b
flabel metal3 1263 8715 1263 8715 0 FreeSans 240 90 0 0 b6a
flabel metal3 1263 10851 1263 10851 0 FreeSans 240 90 0 0 b7a
flabel metal3 1263 10726 1263 10726 0 FreeSans 240 90 0 0 b7b
flabel metal3 1267 12861 1267 12861 0 FreeSans 240 90 0 0 b6a
flabel metal3 1267 12975 1267 12975 0 FreeSans 240 90 0 0 b6b
flabel space 1290 15114 1290 15114 0 FreeSans 240 90 0 0 nca1
flabel space 1292 14993 1292 14993 0 FreeSans 240 90 0 0 ncb1
flabel metal3 1270 17244 1270 17244 0 FreeSans 240 90 0 0 b6a
flabel metal3 1272 17123 1272 17123 0 FreeSans 240 90 0 0 b6b
flabel metal3 1270 19378 1270 19378 0 FreeSans 240 90 0 0 b7b
flabel metal3 1272 19258 1272 19258 0 FreeSans 240 90 0 0 b7a
flabel metal3 1270 21513 1270 21513 0 FreeSans 240 90 0 0 b6b
flabel metal3 1272 21392 1272 21392 0 FreeSans 240 90 0 0 b6a
flabel space 1284 23639 1284 23639 0 FreeSans 240 90 0 0 nca2
flabel space 1286 23518 1286 23518 0 FreeSans 240 90 0 0 ncb2
flabel metal2 6872 30997 7127 31251 0 FreeSans 400 0 0 0 out
port 9 nsew signal output
flabel metal4 s 16541 0 16923 4429 0 FreeSans 1600 270 0 0 dvss
port 14 nsew ground bidirectional
flabel metal4 s 15224 0 15606 4429 0 FreeSans 1600 270 0 0 dvdd
port 13 nsew power bidirectional
flabel metal4 s 792 0 1353 5921 0 FreeSans 1600 270 0 0 avss
port 11 nsew ground bidirectional
flabel metal4 s 792 26880 1429 31244 0 FreeSans 1600 90 0 0 avss
port 11 nsew ground bidirectional
flabel metal4 s 792 5921 1218 26880 0 FreeSans 1600 90 0 0 avss
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16923 31251
<< end >>
