VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rdac3v_8bit
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rdac3v_8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 156.090 BY 84.505 ;
  PIN b0
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 3.475 2.825 3.765 ;
    END
  END b0
  PIN b1
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 11.615 2.825 11.905 ;
    END
  END b1
  PIN b2
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 19.755 2.825 20.045 ;
    END
  END b2
  PIN b3
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 27.895 2.825 28.185 ;
    END
  END b3
  PIN b4
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 36.035 2.825 36.325 ;
    END
  END b4
  PIN b5
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 44.175 2.825 44.465 ;
    END
  END b5
  PIN b6
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 52.315 2.825 52.605 ;
    END
  END b6
  PIN b7
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 60.455 2.825 60.745 ;
    END
  END b7
  PIN out
    ANTENNAGATEAREA 2.400000 ;
    ANTENNADIFFAREA 48.430000 ;
    PORT
      LAYER met2 ;
        RECT 153.635 48.870 156.255 50.145 ;
    END
  END out
  PIN vdd
    ANTENNAGATEAREA 105.000000 ;
    ANTENNADIFFAREA 423.610504 ;
    PORT
      LAYER met4 ;
        RECT -1.000 81.400 18.290 84.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.695 -1.000 34.070 1.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.710 81.400 156.310 84.500 ;
    END
  END vdd
  PIN vss
    ANTENNAGATEAREA 68.250000 ;
    ANTENNADIFFAREA 76.670097 ;
    PORT
      LAYER met4 ;
        RECT -1.000 76.265 26.870 79.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.185 0.330 127.715 2.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.400 77.360 156.290 80.545 ;
    END
  END vss
  PIN ena
    ANTENNAGATEAREA 0.702500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met1 ;
        RECT -1.000 67.695 21.515 67.875 ;
    END
  END ena
  PIN dvdd
    ANTENNADIFFAREA 7.862400 ;
    PORT
      LAYER met2 ;
        RECT -1.000 70.970 2.985 72.695 ;
    END
  END dvdd
  PIN dvss
    ANTENNADIFFAREA 214.649200 ;
    PORT
      LAYER met2 ;
        RECT -1.000 73.455 8.070 75.350 ;
    END
  END dvss
  PIN Vhigh
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER met3 ;
        RECT 34.480 -1.000 35.665 7.215 ;
    END
  END Vhigh
  PIN Vlow
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER met3 ;
        RECT 122.735 -1.000 123.840 7.715 ;
    END
  END Vlow
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 155.600 80.190 ;
      LAYER li1 ;
        RECT 0.330 78.985 156.090 79.960 ;
        RECT 0.330 16.160 156.215 78.985 ;
        RECT 0.330 0.430 156.090 16.160 ;
      LAYER met1 ;
        RECT 0.330 78.985 156.090 79.970 ;
        RECT 0.330 68.155 156.215 78.985 ;
        RECT 21.795 67.415 156.215 68.155 ;
        RECT 0.330 61.025 156.215 67.415 ;
        RECT 3.105 60.175 156.215 61.025 ;
        RECT 0.330 52.885 156.215 60.175 ;
        RECT 3.105 52.035 156.215 52.885 ;
        RECT 0.330 44.745 156.215 52.035 ;
        RECT 3.105 43.895 156.215 44.745 ;
        RECT 0.330 36.605 156.215 43.895 ;
        RECT 3.105 35.755 156.215 36.605 ;
        RECT 0.330 28.465 156.215 35.755 ;
        RECT 3.105 27.615 156.215 28.465 ;
        RECT 0.330 20.325 156.215 27.615 ;
        RECT 3.105 19.475 156.215 20.325 ;
        RECT 0.330 16.160 156.215 19.475 ;
        RECT 0.330 12.185 156.090 16.160 ;
        RECT 3.105 11.335 156.090 12.185 ;
        RECT 0.330 4.045 156.090 11.335 ;
        RECT 3.105 3.195 156.090 4.045 ;
        RECT 0.330 0.000 156.090 3.195 ;
        RECT 131.370 -0.110 135.250 0.000 ;
      LAYER met2 ;
        RECT 1.520 75.630 155.980 84.505 ;
        RECT 8.350 73.175 155.980 75.630 ;
        RECT 1.520 72.975 155.980 73.175 ;
        RECT 3.265 70.690 155.980 72.975 ;
        RECT 1.520 50.425 155.980 70.690 ;
        RECT 1.520 48.590 153.355 50.425 ;
        RECT 1.520 0.000 155.980 48.590 ;
        RECT 7.160 -0.110 135.250 0.000 ;
      LAYER met3 ;
        RECT 4.130 8.115 155.980 84.505 ;
        RECT 4.130 7.615 122.335 8.115 ;
        RECT 4.130 1.550 34.080 7.615 ;
        RECT 4.130 0.000 31.295 1.550 ;
        RECT 36.065 0.000 122.335 7.615 ;
        RECT 124.240 2.680 155.980 8.115 ;
        RECT 124.185 -1.000 125.985 0.330 ;
        RECT 128.115 0.000 155.980 2.680 ;
      LAYER met4 ;
        RECT 18.690 81.000 138.310 84.500 ;
        RECT 18.160 80.945 156.090 81.000 ;
        RECT 18.160 80.035 134.000 80.945 ;
        RECT 27.270 76.960 134.000 80.035 ;
        RECT 156.290 78.415 156.305 80.545 ;
        RECT 27.270 75.865 156.090 76.960 ;
        RECT 18.160 0.330 156.090 75.865 ;
      LAYER met5 ;
        RECT 38.415 8.850 114.635 70.550 ;
  END
END sky130_ef_ip__rdac3v_8bit
END LIBRARY

