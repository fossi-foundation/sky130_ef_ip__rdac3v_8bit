VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rdac3v_8bit
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rdac3v_8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 84.615 BY 156.255 ;
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 80.740 0.000 81.030 0.910 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 72.600 0.000 72.890 0.910 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 64.460 0.000 64.750 0.910 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 56.320 0.000 56.610 0.910 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 48.180 0.000 48.470 0.910 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 40.040 0.000 40.330 0.910 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 31.900 0.000 32.190 0.910 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 23.760 0.000 24.050 0.910 ;
    END
  END b[7]
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.400000 ;
    ANTENNADIFFAREA 48.430000 ;
    PORT
      LAYER met2 ;
        RECT 34.360 153.635 35.635 156.255 ;
    END
  END out
  PIN avdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.005 0.000 3.105 156.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.495 31.695 84.615 34.070 ;
    END
  END avdd
  PIN avss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 82.225 124.185 84.615 125.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.960 0.000 6.765 29.605 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.960 134.400 7.145 156.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.960 29.605 6.090 134.400 ;
    END
  END avss
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.702500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 16.630 0.000 16.810 0.920 ;
    END
  END ena
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 11.810 0.000 13.535 2.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.120 0.000 78.030 22.145 ;
    END
  END dvdd
  PIN dvss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 9.155 0.000 11.050 8.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.705 0.000 84.615 22.145 ;
    END
  END dvss
  PIN Vhigh
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER met3 ;
        RECT 77.290 34.480 84.615 35.665 ;
    END
  END Vhigh
  PIN Vlow
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER met3 ;
        RECT 76.790 122.735 84.615 123.840 ;
    END
  END Vlow
  OBS
      LAYER nwell ;
        RECT 4.315 0.000 84.505 156.060 ;
      LAYER li1 ;
        RECT 4.990 156.255 68.345 156.675 ;
        RECT 4.545 0.330 84.075 156.255 ;
      LAYER met1 ;
        RECT 4.990 156.255 68.345 156.675 ;
        RECT 4.535 0.330 84.615 156.255 ;
      LAYER met2 ;
        RECT 0.000 153.355 34.080 155.980 ;
        RECT 35.915 153.355 84.615 155.980 ;
        RECT 0.000 8.350 84.615 153.355 ;
        RECT 0.000 0.610 8.875 8.350 ;
        RECT 11.330 3.265 84.615 8.350 ;
        RECT 11.330 0.610 11.530 3.265 ;
        RECT 13.815 1.200 84.615 3.265 ;
        RECT 13.815 0.610 16.350 1.200 ;
        RECT 17.090 1.190 84.615 1.200 ;
        RECT 17.090 0.610 23.480 1.190 ;
        RECT 24.330 0.610 31.620 1.190 ;
        RECT 32.470 0.610 39.760 1.190 ;
        RECT 40.610 0.610 47.900 1.190 ;
        RECT 48.750 0.610 56.040 1.190 ;
        RECT 56.890 0.610 64.180 1.190 ;
        RECT 65.030 0.610 72.320 1.190 ;
        RECT 73.170 0.610 80.460 1.190 ;
        RECT 81.310 0.610 84.615 1.190 ;
      LAYER met3 ;
        RECT 0.000 126.385 84.610 155.980 ;
        RECT 0.000 124.240 81.825 126.385 ;
        RECT 0.000 122.335 76.390 124.240 ;
        RECT 0.000 36.065 84.610 122.335 ;
        RECT 0.000 34.080 76.890 36.065 ;
        RECT 0.000 31.295 81.095 34.080 ;
        RECT 0.000 0.610 84.610 31.295 ;
      LAYER met4 ;
        RECT 7.545 134.000 84.175 136.810 ;
        RECT 6.490 30.005 84.175 134.000 ;
        RECT 7.165 22.545 84.175 30.005 ;
        RECT 7.165 18.160 75.720 22.545 ;
        RECT 78.430 18.160 82.305 22.545 ;
      LAYER met5 ;
        RECT 13.955 38.415 75.655 114.635 ;
  END
END sky130_ef_ip__rdac3v_8bit
END LIBRARY

